module A;
always_comb begin
    case (x)
        1: y = 0;
    endcase

end
always_ff begin
    case (x)
        1: y = 0;
    endcase
end
endmodule
